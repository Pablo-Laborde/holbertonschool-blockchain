HBLK0.3              ��[                                               Holberton School�,&ȵF9c]��*�ԍ� 	�����/QX����       %�g            �,&ȵF9c]��*�ԍ� 	�����/QX   Node 1�ȉ�!W鶰����Hټ�N'��9F���"k9O   >�8����	�f,�#'Y,wHf����CA�                                                                                                                                                                              2   �t{������q<���_����&}����J��HU�l��/���@ˋ������ᝫ�q�`9G�֙`��9�&��o�Gl�Y����T!�       %�g            �ȉ�!W鶰����Hټ�N'��9F���"k9O   Node 2aK��B���F1���ws�#j�vӋ��� =E�d   �f��0�Ec6b��]:kWy����Í腯F���                                                                                                                                                                              2   ��n+y��A�Qz 4T�*j�eBk.��4�`�(�#nI�)��[����KG��h. �K�2W^y��C 2׾Æ>;�&��d� ~�"       %�g            aK��B���F1���ws�#j�vӋ��� =E�d   Node 3�C��M�Ћ�`l�i��G9���}Cj %]   9qdT��8>�ll4���.G�m��5�CI��p��V                                                                                                                                                                              2   ����3Ϫ�_;~�鏝@!WǮ��
�,��>�=+��sn*[��M�W'�4��N�u�[� eք��˝�zP��6	�
�L�}(ش |�s���=       %�g            �C��M�Ћ�`l�i��G9���}Cj %]   Node 4�4>n�e���?RS����c���^�߳*${�   �@�V��n��&��*�h ���M���ii��                                                                                                                                                                              2   lG�L��6Q�ܩP�������wB��L0��mn�q��8:�uE
'��o}�M� ���&�~�l��\�r��Q)9[}��=��C�7���bPi�/e�|P       %�g            �4>n�e���?RS����c���^�߳*${�   Node 5�#}-�8q"͔i�i�"�TZ�}�nE ��$   ���R*t/���PO���<pn�㙨�����%��                                                                                                                                                                              2   ���f��<�Dݡ���GC�H���V��<�NY�,俔�It�&�d%>_�/�������4q��4�R�$(�F�0�n�dK/�v�Wu�KK��      %�g           �#}-�8q"͔i�i�"�TZ�}�nE ��$   Node 6]|�_��:FSJ�7��LSU�$\��������   ;c>����z�ʢ6�20֌EIi����'(�;�                                                                                                                                                                              2   /R��aQ7=������`���(���@U���=x���>zI�[zշ����"����z�(5g+Ot��Áݕ�h�ol՘W���Y`�;/�py۰C�=�ȉ�!W鶰����Hټ�N'��9F���"k9O>�8����	�f,�#'Y,wHf����CA�2   �t{������q<���_����&}����J��HU�l��/���@ˋ������ᝫ�q�`9G�֙`��9�&��o�Gl�Y����T!�aK��B���F1���ws�#j�vӋ��� =E�d�f��0�Ec6b��]:kWy����Í腯F���2   ��n+y��A�Qz 4T�*j�eBk.��4�`�(�#nI�)��[����KG��h. �K�2W^y��C 2׾Æ>;�&��d� ~�"�C��M�Ћ�`l�i��G9���}Cj %]9qdT��8>�ll4���.G�m��5�CI��p��V2   ����3Ϫ�_;~�鏝@!WǮ��
�,��>�=+��sn*[��M�W'�4��N�u�[� eք��˝�zP��6	�
�L�}(ش |�s���=�4>n�e���?RS����c���^�߳*${�@�V��n��&��*�h ���M���ii��2   lG�L��6Q�ܩP�������wB��L0��mn�q��8:�uE
'��o}�M� ���&�~�l��\�r��Q)9[}��=��C�7���bPi�/e�|P�#}-�8q"͔i�i�"�TZ�}�nE ��$���R*t/���PO���<pn�㙨�����%��2   ���f��<�Dݡ���GC�H���V��<�NY�,俔�It�&�d%>_�/�������4q��4�R�$(�F�0�n�dK/�v�Wu�KK��]|�_��:FSJ�7��LSU�$\��������;c>����z�ʢ6�20֌EIi����'(�;�2   /R��aQ7=������`���(���@U���=x���>zI�[zշ����"����z�(5g+Ot��Áݕ�h�ol՘W���Y`�;/�py۰C�=