HBLK0.3              ��[                                               Holberton School�,&ȵF9c]��*�ԍ� 	�����/QX����       ��g            �,&ȵF9c]��*�ԍ� 	�����/QX   Node 1�O�l)=���<��C&P�J���DI_o'�[��k   ����G��`���I/ޣH���k��uy^��5                                                                                                                                                                              2   Pd���;*��9p������|���5�QC5lb�����L�Wpd�+G��:2�"�M��O�������j?A�.�+�"H�F��)��Q�p4
       ��g            �O�l)=���<��C&P�J���DI_o'�[��k   Node 2rr�p {����{���1_^&=Z�:��C/�K   �w����[���"�!��q�~_��WY��@��V                                                                                                                                                                              2   ���i�q5������[�K�0�&z��2���B��b^@~�6W[Ȉa��a��N?�z��x�A��\�D�y����L���B;�������mv-       ��g            rr�p {����{���1_^&=Z�:��C/�K   Node 3�9��7?�� �����<t۷^��*xN   �T�����\�>U`>7駙�}�
w�$�[��                                                                                                                                                                              2   ��u/��L��Q�m����/����5@��� �ƏP�+A ��+.j���w~U���J�^y�m��פ��E�7��8�m�#�k��/j       ��g            �9��7?�� �����<t۷^��*xN   Node 4�f\�F��5;�v��-��1�疶/��Mo��\�I1   �V��m���;`���b6/1t���$	��6�*b^                                                                                                                                                                              2   '3���~L��o�2y�}�^�zꠚ�����xo)|�q�9\'����^w&�T��D,`@�M��|�S'Q>����0��_(�-��``yl��~       ��g            �f\�F��5;�v��-��1�疶/��Mo��\�I1   Node 5{�����F����Z�����l�,�N   �z�����3�#[�.]��Î�{*`��;��t�                                                                                                                                                                              2   J�w��n`�|�� ���>��C@5���PY��`�ݨ�2ze���m��,Ӛ����HEb�-�<#M����n_�:Ԃ��l�4O�޲E�>      ��g            {�����F����Z�����l�,�N   Node 6^��D��R�S�����xIj�r3�"��   �l_�~�(t�Z~{���W�}{�!�=2�Q;E�B                                                                                                                                                                              2   N��v��Q�w���'���L�C�_e��a�tTp�������밁{Ns\6�QS�xϏ�S�I�T��2��{�|����w�����ij��W�|�O�l)=���<��C&P�J���DI_o'�[��k����G��`���I/ޣH���k��uy^��52   Pd���;*��9p������|���5�QC5lb�����L�Wpd�+G��:2�"�M��O�������j?A�.�+�"H�F��)��Q�p4
rr�p {����{���1_^&=Z�:��C/�K�w����[���"�!��q�~_��WY��@��V2   ���i�q5������[�K�0�&z��2���B��b^@~�6W[Ȉa��a��N?�z��x�A��\�D�y����L���B;�������mv-�9��7?�� �����<t۷^��*xN�T�����\�>U`>7駙�}�
w�$�[��2   ��u/��L��Q�m����/����5@��� �ƏP�+A ��+.j���w~U���J�^y�m��פ��E�7��8�m�#�k��/j�f\�F��5;�v��-��1�疶/��Mo��\�I1�V��m���;`���b6/1t���$	��6�*b^2   '3���~L��o�2y�}�^�zꠚ�����xo)|�q�9\'����^w&�T��D,`@�M��|�S'Q>����0��_(�-��``yl��~{�����F����Z�����l�,�N�z�����3�#[�.]��Î�{*`��;��t�2   J�w��n`�|�� ���>��C@5���PY��`�ݨ�2ze���m��,Ӛ����HEb�-�<#M����n_�:Ԃ��l�4O�޲E�>^��D��R�S�����xIj�r3�"���l_�~�(t�Z~{���W�}{�!�=2�Q;E�B2   N��v��Q�w���'���L�C�_e��a�tTp�������밁{Ns\6�QS�xϏ�S�I�T��2��{�|����w�����ij��W�|